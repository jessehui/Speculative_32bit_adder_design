-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition
-- Created on Wed Apr 27 12:26:06 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY judge_fsm IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        co : IN STD_LOGIC := '0';
        mi : OUT STD_LOGIC;
        ctl_reg : OUT STD_LOGIC
    );
END judge_fsm;

ARCHITECTURE BEHAVIOR OF judge_fsm IS
    TYPE type_fstate IS (A,B,C);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,co)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            mi <= '0';
            ctl_reg <= '0';
        ELSE
            mi <= '0';
            ctl_reg <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((co = '1')) THEN
                        reg_fstate <= C;
                    ELSIF ((co = '0')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    ctl_reg <= '1';

                    mi <= '0';
                WHEN B =>
                    IF ((co = '0')) THEN
                        reg_fstate <= A;
                    ELSIF ((co = '1')) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B;
                    END IF;

                    ctl_reg <= '0';

                    mi <= '0';
                WHEN C =>
                    IF ((co = '0')) THEN
                        reg_fstate <= B;
                    ELSIF ((co = '1')) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    ctl_reg <= '1';

                    mi <= '1';
                WHEN OTHERS => 
                    mi <= 'X';
                    ctl_reg <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
